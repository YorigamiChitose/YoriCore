/* verilator lint_off NULLPORT */
module SimInfo (
  input       clock,
  input       reset,
  input       SI_PC_IF_ioValid,
  input       SI_IF_ID_ioValid,
  input       SI_ID_EX_ioValid,
  input       SI_EX_WB_ioValid,
  input [3:0] SI_EX_WB_excType
);

endmodule
/* verilator lint_on NULLPORT */